`ifndef IMMEDIATE_SVH
`define IMMEDIATE_SVH

typedef enum logic [2:0] {
  IMM_I,
  IMM_S,
  IMM_B,
  IMM_U,
  IMM_J
} immediate_e;

`endif
