`ifndef INSTRUCTIONS_VH
`define INSTRUCTIONS_VH

localparam unsigned INSTRUCTION_NOP = 32'h00000013;

`endif
