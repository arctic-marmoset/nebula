package addressing;

  localparam bit [31:0] BaseAddress = 'h80000000;

endpackage
