package types;

  typedef logic [63:0] dword_t;
  typedef logic [31:0] word_t;
  typedef logic [15:0] hword_t;

  typedef word_t x_t;

endpackage
