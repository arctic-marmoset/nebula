`ifndef WRITEBACK_SVH
`define WRITEBACK_SVH

typedef enum logic [0:0] {
    WB_SRC_ALU,
    WB_SRC_PC_NEXT_SEQUENTIAL
} writeback_source_e;

`endif
