`ifndef INSTRUCTIONS_VH
`define INSTRUCTIONS_VH

/* verilator lint_off UNUSEDPARAM */
localparam logic [31:0] INSTRUCTION_NOP = 32'h00000013;
localparam logic [31:0] INSTRUCTION_WFI = 32'h10500073;
/* verilator lint_on UNUSEDPARAM */

`endif
